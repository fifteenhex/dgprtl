module fontrom
(
    input logic clk,
    input logic [11:0] addr,
    output logic [7:0] data
);

    reg [31:8] data_discard;
    reg [7:0] rom_data;

    pROM bram_prom_0 (
        .DO({data_discard, data}),
        .CLK(clk),
        .OCE('1),
        .CE('1),
        .RESET('0),
        .AD({addr[10:0],3'b000})
    );
    defparam bram_prom_0.READ_MODE=1'b0;
    defparam bram_prom_0.BIT_WIDTH = 8;
    defparam bram_prom_0.RESET_MODE="ASYNC";

defparam bram_prom_0.INIT_RAM_00=256'h000000007e818199bd8181a5817e000000000000000000000000000000000000;
defparam bram_prom_0.INIT_RAM_01=256'h0000000010387cfefefefe6c00000000000000007effffe7c3ffffdbff7e0000;
defparam bram_prom_0.INIT_RAM_02=256'h000000003c1818e7e7e73c3c18000000000000000010387cfe7c381000000000;
defparam bram_prom_0.INIT_RAM_03=256'h000000000000183c3c18000000000000000000003c18187effff7e3c18000000;
defparam bram_prom_0.INIT_RAM_04=256'h00000000003c664242663c0000000000ffffffffffffe7c3c3e7ffffffffffff;
defparam bram_prom_0.INIT_RAM_05=256'h0000000078cccccccc78321a0e1e0000ffffffffffc399bdbd99c3ffffffffff;
defparam bram_prom_0.INIT_RAM_06=256'h00000000e0f070303030303f333f00000000000018187e183c666666663c0000;
defparam bram_prom_0.INIT_RAM_07=256'h000000001818db3ce73cdb1818000000000000c0e6e767636363637f637f0000;
defparam bram_prom_0.INIT_RAM_08=256'h0000000002060e1e3efe3e1e0e0602000000000080c0e0f0f8fef8f0e0c08000;
defparam bram_prom_0.INIT_RAM_09=256'h000000006666006666666666666600000000000000183c7e1818187e3c180000;
defparam bram_prom_0.INIT_RAM_0A=256'h0000007cc60c386cc6c66c3860c67c00000000001b1b1b1b1b7bdbdbdb7f0000;
defparam bram_prom_0.INIT_RAM_0B=256'h000000007e183c7e1818187e3c18000000000000fefefefe0000000000000000;
defparam bram_prom_0.INIT_RAM_0C=256'h00000000183c7e18181818181818000000000000181818181818187e3c180000;
defparam bram_prom_0.INIT_RAM_0D=256'h0000000000003060fe60300000000000000000000000180cfe0c180000000000;
defparam bram_prom_0.INIT_RAM_0E=256'h0000000000002466ff66240000000000000000000000fec0c0c0000000000000;
defparam bram_prom_0.INIT_RAM_0F=256'h00000000001038387c7cfefe000000000000000000fefe7c7c38381000000000;
defparam bram_prom_0.INIT_RAM_10=256'h000000001818001818183c3c3c18000000000000000000000000000000000000;
defparam bram_prom_0.INIT_RAM_11=256'h000000006c6cfe6c6c6cfe6c6c00000000000000000000000000002466666600;
defparam bram_prom_0.INIT_RAM_12=256'h0000000086c66030180cc6c200000000000018187cc68606067cc0c2c67c1818;
defparam bram_prom_0.INIT_RAM_13=256'h000000000000000000000060303030000000000076ccccccdc76386c6c380000;
defparam bram_prom_0.INIT_RAM_14=256'h0000000030180c0c0c0c0c0c18300000000000000c18303030303030180c0000;
defparam bram_prom_0.INIT_RAM_15=256'h00000000000018187e18180000000000000000000000663cff3c660000000000;
defparam bram_prom_0.INIT_RAM_16=256'h0000000000000000fe0000000000000000000030181818000000000000000000;
defparam bram_prom_0.INIT_RAM_17=256'h0000000080c06030180c06020000000000000000181800000000000000000000;
defparam bram_prom_0.INIT_RAM_18=256'h000000007e1818181818187838180000000000003c66c3c3dbdbc3c3663c0000;
defparam bram_prom_0.INIT_RAM_19=256'h000000007cc60606063c0606c67c000000000000fec6c06030180c06c67c0000;
defparam bram_prom_0.INIT_RAM_1A=256'h000000007cc6060606fcc0c0c0fe0000000000001e0c0c0cfecc6c3c1c0c0000;
defparam bram_prom_0.INIT_RAM_1B=256'h0000000030303030180c0606c6fe0000000000007cc6c6c6c6fcc0c060380000;
defparam bram_prom_0.INIT_RAM_1C=256'h00000000780c0606067ec6c6c67c0000000000007cc6c6c6c67cc6c6c67c0000;
defparam bram_prom_0.INIT_RAM_1D=256'h0000000030181800000018180000000000000000001818000000181800000000;
defparam bram_prom_0.INIT_RAM_1E=256'h000000000000007e00007e000000000000000000060c18306030180c06000000;
defparam bram_prom_0.INIT_RAM_1F=256'h000000001818001818180cc6c67c0000000000006030180c060c183060000000;
defparam bram_prom_0.INIT_RAM_20=256'h00000000c6c6c6c6fec6c66c38100000000000007cc0dcdededec6c67c000000;
defparam bram_prom_0.INIT_RAM_21=256'h000000003c66c2c0c0c0c0c2663c000000000000fc666666667c666666fc0000;
defparam bram_prom_0.INIT_RAM_22=256'h00000000fe6662606878686266fe000000000000f86c6666666666666cf80000;
defparam bram_prom_0.INIT_RAM_23=256'h000000003a66c6c6dec0c0c2663c000000000000f06060606878686266fe0000;
defparam bram_prom_0.INIT_RAM_24=256'h000000003c18181818181818183c000000000000c6c6c6c6c6fec6c6c6c60000;
defparam bram_prom_0.INIT_RAM_25=256'h00000000e666666c78786c6666e600000000000078cccccc0c0c0c0c0c1e0000;
defparam bram_prom_0.INIT_RAM_26=256'h00000000c3c3c3c3c3dbffffe7c3000000000000fe6662606060606060f00000;
defparam bram_prom_0.INIT_RAM_27=256'h000000007cc6c6c6c6c6c6c6c67c000000000000c6c6c6c6cedefef6e6c60000;
defparam bram_prom_0.INIT_RAM_28=256'h00000e0c7cded6c6c6c6c6c6c67c000000000000f0606060607c666666fc0000;
defparam bram_prom_0.INIT_RAM_29=256'h000000007cc6c6060c3860c6c67c000000000000e66666666c7c666666fc0000;
defparam bram_prom_0.INIT_RAM_2A=256'h000000007cc6c6c6c6c6c6c6c6c60000000000003c18181818181899dbff0000;
defparam bram_prom_0.INIT_RAM_2B=256'h000000006666ffdbdbc3c3c3c3c3000000000000183c66c3c3c3c3c3c3c30000;
defparam bram_prom_0.INIT_RAM_2C=256'h000000003c181818183c66c3c3c3000000000000c3c3663c18183c66c3c30000;
defparam bram_prom_0.INIT_RAM_2D=256'h000000003c30303030303030303c000000000000ffc3c16030180c86c3ff0000;
defparam bram_prom_0.INIT_RAM_2E=256'h000000003c0c0c0c0c0c0c0c0c3c00000000000002060e1c3870e0c080000000;
defparam bram_prom_0.INIT_RAM_2F=256'h0000ff00000000000000000000000000000000000000000000000000c66c3810;
defparam bram_prom_0.INIT_RAM_30=256'h0000000076cccccc7c0c78000000000000000000000000000000000000183030;
defparam bram_prom_0.INIT_RAM_31=256'h000000007cc6c0c0c0c67c0000000000000000007c666666666c786060e00000;
defparam bram_prom_0.INIT_RAM_32=256'h000000007cc6c0c0fec67c00000000000000000076cccccccc6c3c0c0c1c0000;
defparam bram_prom_0.INIT_RAM_33=256'h0078cc0c7ccccccccccc76000000000000000000f060606060f060646c380000;
defparam bram_prom_0.INIT_RAM_34=256'h000000003c181818181838001818000000000000e666666666766c6060e00000;
defparam bram_prom_0.INIT_RAM_35=256'h00000000e6666c78786c666060e00000003c66660606060606060e0006060000;
defparam bram_prom_0.INIT_RAM_36=256'h00000000dbdbdbdbdbffe60000000000000000003c1818181818181818380000;
defparam bram_prom_0.INIT_RAM_37=256'h000000007cc6c6c6c6c67c000000000000000000666666666666dc0000000000;
defparam bram_prom_0.INIT_RAM_38=256'h001e0c0c7ccccccccccc76000000000000f060607c6666666666dc0000000000;
defparam bram_prom_0.INIT_RAM_39=256'h000000007cc60c3860c67c000000000000000000f06060606676dc0000000000;
defparam bram_prom_0.INIT_RAM_3A=256'h0000000076cccccccccccc0000000000000000001c3630303030fc3030100000;
defparam bram_prom_0.INIT_RAM_3B=256'h0000000066ffdbdbc3c3c3000000000000000000183c66c3c3c3c30000000000;
defparam bram_prom_0.INIT_RAM_3C=256'h00f80c067ec6c6c6c6c6c6000000000000000000c3663c183c66c30000000000;
defparam bram_prom_0.INIT_RAM_3D=256'h000000000e18181818701818180e000000000000fec6603018ccfe0000000000;
defparam bram_prom_0.INIT_RAM_3E=256'h0000000070181818180e18181870000000000000181818181800181818180000;
defparam bram_prom_0.INIT_RAM_3F=256'h0000000000fec6c6c66c381000000000000000000000000000000000dc760000;

endmodule
